@00000000
8C 08 04 00 8C 0A 02 00 00 00 00 00 11 0A 00 06 
00 00 00 00 8C 09 08 00 00 00 00 00 AC 09 04 00 
08 00 00 00 AC 09 08 00 8C 08 02 01 31 4A 00 00 
21 08 FF FF 11 0A 00 03 00 00 00 00 08 00 00 0C 
00 00 00 00 8C 08 02 02 8C 0A 02 11 8D 09 00 00 
00 00 00 00 AC 09 04 00 21 08 00 01 11 0A FF E8 
00 00 00 00 08 00 00 13 00 00 00 00 08 00 00 00 
00 00 00 00 
@00400098
00 00 01 00 01 01 00 01 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 

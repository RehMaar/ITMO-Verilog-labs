@00000200
00 00 00 01 00 0F 42 40 48 65 6C 6C 6F 2C 20 77 
6F 72 6C 64 21 0A 0D 
@00400098
00 00 01 00 01 01 00 01 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 

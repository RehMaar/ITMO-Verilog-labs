@00000200
00 00 00 01 00 00 01 00 00 00 00 48 00 00 00 65 
00 00 00 6C 00 00 00 6C 00 00 00 6F 00 00 00 2C 
00 00 00 20 00 00 00 77 00 00 00 6F 00 00 00 72 
00 00 00 6C 00 00 00 64 00 00 00 21 00 00 00 0D 
00 00 00 0A 
@00400098
00 00 01 00 01 01 00 01 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 

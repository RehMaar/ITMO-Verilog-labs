@00000000
8C 08 02 00 00 00 00 00 01 28 48 24 AC 09 04 00 
8C 08 02 01 00 00 00 00 01 48 50 24 AC 0A 04 00 
8C 08 02 02 00 00 00 00 01 28 48 24 AC 09 04 00 
01 48 50 24 AC 0A 04 00 8C 08 02 03 00 00 00 00 
01 28 48 24 AC 09 04 00 01 48 50 24 AC 0A 04 00 
@00400098
00 00 01 00 01 01 00 01 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 

@00000200
00 01 00 01 11 01 11 11 00 00 00 00 11 11 11 11 
@00400098
00 00 01 00 01 01 00 01 00 00 00 00 00 00 00 00 
00 00 00 00 00 00 00 00 
